module OneHotDecoder_1(
  input  [2:0] io_in,
  output [7:0] io_out
);
  wire  bools_0; // @[OneHotDecoder.scala 14:46]
  wire  bools_1; // @[OneHotDecoder.scala 14:46]
  wire  bools_2; // @[OneHotDecoder.scala 14:46]
  wire  bools_3; // @[OneHotDecoder.scala 14:46]
  wire  bools_4; // @[OneHotDecoder.scala 14:46]
  wire  bools_5; // @[OneHotDecoder.scala 14:46]
  wire  bools_6; // @[OneHotDecoder.scala 14:46]
  wire  bools_7; // @[OneHotDecoder.scala 14:46]
  wire [3:0] _T_40; // @[OneHotDecoder.scala 16:25]
  wire [3:0] _T_43; // @[OneHotDecoder.scala 16:25]
  assign bools_0 = io_in == 3'h0; // @[OneHotDecoder.scala 14:46]
  assign bools_1 = io_in == 3'h1; // @[OneHotDecoder.scala 14:46]
  assign bools_2 = io_in == 3'h2; // @[OneHotDecoder.scala 14:46]
  assign bools_3 = io_in == 3'h3; // @[OneHotDecoder.scala 14:46]
  assign bools_4 = io_in == 3'h4; // @[OneHotDecoder.scala 14:46]
  assign bools_5 = io_in == 3'h5; // @[OneHotDecoder.scala 14:46]
  assign bools_6 = io_in == 3'h6; // @[OneHotDecoder.scala 14:46]
  assign bools_7 = io_in == 3'h7; // @[OneHotDecoder.scala 14:46]
  assign _T_40 = {bools_3,bools_2,bools_1,bools_0}; // @[OneHotDecoder.scala 16:25]
  assign _T_43 = {bools_7,bools_6,bools_5,bools_4}; // @[OneHotDecoder.scala 16:25]
  assign io_out = {_T_43,_T_40}; // @[OneHotDecoder.scala 16:10]
endmodule
module OneHotEncoder(
  input        io_in_1,
  input        io_in_2,
  input        io_in_3,
  input        io_in_4,
  input        io_in_5,
  input        io_in_6,
  input        io_in_7,
  input        io_in_8,
  input        io_in_9,
  input        io_in_10,
  input        io_in_11,
  input        io_in_12,
  input        io_in_13,
  input        io_in_14,
  output [3:0] io_out
);
  wire [3:0] _T_74; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_76; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_89; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_91; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_104; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_106; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_119; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_121; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_134; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_136; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_149; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_151; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_164; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_166; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_179; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_181; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_194; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_196; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_209; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_211; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_224; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_226; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_239; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_241; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_254; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_256; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_269; // @[OneHotEncoder.scala 12:94]
  wire [3:0] _T_271; // @[OneHotEncoder.scala 12:97]
  wire [3:0] _T_273; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_274; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_275; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_276; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_277; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_278; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_279; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_280; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_281; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_282; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_283; // @[OneHotEncoder.scala 12:113]
  wire [3:0] _T_284; // @[OneHotEncoder.scala 12:113]
  assign _T_74 = {io_in_1,io_in_1,io_in_1,io_in_1}; // @[OneHotEncoder.scala 12:94]
  assign _T_76 = _T_74 & 4'h1; // @[OneHotEncoder.scala 12:97]
  assign _T_89 = {io_in_2,io_in_2,io_in_2,io_in_2}; // @[OneHotEncoder.scala 12:94]
  assign _T_91 = _T_89 & 4'h2; // @[OneHotEncoder.scala 12:97]
  assign _T_104 = {io_in_3,io_in_3,io_in_3,io_in_3}; // @[OneHotEncoder.scala 12:94]
  assign _T_106 = _T_104 & 4'h3; // @[OneHotEncoder.scala 12:97]
  assign _T_119 = {io_in_4,io_in_4,io_in_4,io_in_4}; // @[OneHotEncoder.scala 12:94]
  assign _T_121 = _T_119 & 4'h4; // @[OneHotEncoder.scala 12:97]
  assign _T_134 = {io_in_5,io_in_5,io_in_5,io_in_5}; // @[OneHotEncoder.scala 12:94]
  assign _T_136 = _T_134 & 4'h5; // @[OneHotEncoder.scala 12:97]
  assign _T_149 = {io_in_6,io_in_6,io_in_6,io_in_6}; // @[OneHotEncoder.scala 12:94]
  assign _T_151 = _T_149 & 4'h6; // @[OneHotEncoder.scala 12:97]
  assign _T_164 = {io_in_7,io_in_7,io_in_7,io_in_7}; // @[OneHotEncoder.scala 12:94]
  assign _T_166 = _T_164 & 4'h7; // @[OneHotEncoder.scala 12:97]
  assign _T_179 = {io_in_8,io_in_8,io_in_8,io_in_8}; // @[OneHotEncoder.scala 12:94]
  assign _T_181 = _T_179 & 4'h8; // @[OneHotEncoder.scala 12:97]
  assign _T_194 = {io_in_9,io_in_9,io_in_9,io_in_9}; // @[OneHotEncoder.scala 12:94]
  assign _T_196 = _T_194 & 4'h9; // @[OneHotEncoder.scala 12:97]
  assign _T_209 = {io_in_10,io_in_10,io_in_10,io_in_10}; // @[OneHotEncoder.scala 12:94]
  assign _T_211 = _T_209 & 4'ha; // @[OneHotEncoder.scala 12:97]
  assign _T_224 = {io_in_11,io_in_11,io_in_11,io_in_11}; // @[OneHotEncoder.scala 12:94]
  assign _T_226 = _T_224 & 4'hb; // @[OneHotEncoder.scala 12:97]
  assign _T_239 = {io_in_12,io_in_12,io_in_12,io_in_12}; // @[OneHotEncoder.scala 12:94]
  assign _T_241 = _T_239 & 4'hc; // @[OneHotEncoder.scala 12:97]
  assign _T_254 = {io_in_13,io_in_13,io_in_13,io_in_13}; // @[OneHotEncoder.scala 12:94]
  assign _T_256 = _T_254 & 4'hd; // @[OneHotEncoder.scala 12:97]
  assign _T_269 = {io_in_14,io_in_14,io_in_14,io_in_14}; // @[OneHotEncoder.scala 12:94]
  assign _T_271 = _T_269 & 4'he; // @[OneHotEncoder.scala 12:97]
  assign _T_273 = _T_76 | _T_91; // @[OneHotEncoder.scala 12:113]
  assign _T_274 = _T_273 | _T_106; // @[OneHotEncoder.scala 12:113]
  assign _T_275 = _T_274 | _T_121; // @[OneHotEncoder.scala 12:113]
  assign _T_276 = _T_275 | _T_136; // @[OneHotEncoder.scala 12:113]
  assign _T_277 = _T_276 | _T_151; // @[OneHotEncoder.scala 12:113]
  assign _T_278 = _T_277 | _T_166; // @[OneHotEncoder.scala 12:113]
  assign _T_279 = _T_278 | _T_181; // @[OneHotEncoder.scala 12:113]
  assign _T_280 = _T_279 | _T_196; // @[OneHotEncoder.scala 12:113]
  assign _T_281 = _T_280 | _T_211; // @[OneHotEncoder.scala 12:113]
  assign _T_282 = _T_281 | _T_226; // @[OneHotEncoder.scala 12:113]
  assign _T_283 = _T_282 | _T_241; // @[OneHotEncoder.scala 12:113]
  assign _T_284 = _T_283 | _T_256; // @[OneHotEncoder.scala 12:113]
  assign io_out = _T_284 | _T_271; // @[OneHotEncoder.scala 12:10]
endmodule
module InstDecoder(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  output [3:0]  io_aluOPCode,
  output [4:0]  io_regInfos_0_regIdx,
  output        io_regInfos_0_need,
  output [4:0]  io_regInfos_1_regIdx,
  output        io_regInfos_1_need,
  output [4:0]  io_regInfos_2_regIdx,
  output        io_regInfos_2_need,
  output [4:0]  io_regInfos_3_regIdx,
  output        io_regInfos_3_need
);
  wire [2:0] decoder_3_8_io_in; // @[InstDecoder.scala 41:27]
  wire [7:0] decoder_3_8_io_out; // @[InstDecoder.scala 41:27]
  wire  alu_op_encoder_io_in_1; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_2; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_3; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_4; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_5; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_6; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_7; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_8; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_9; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_10; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_11; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_12; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_13; // @[InstDecoder.scala 288:30]
  wire  alu_op_encoder_io_in_14; // @[InstDecoder.scala 288:30]
  wire [3:0] alu_op_encoder_io_out; // @[InstDecoder.scala 288:30]
  wire [6:0] _T_37; // @[InstDecoder.scala 69:38]
  wire  func7_op_0; // @[InstDecoder.scala 69:46]
  wire  func7_op_100000; // @[InstDecoder.scala 70:46]
  wire [5:0] _T_41; // @[InstDecoder.scala 71:38]
  wire  func6_op_0; // @[InstDecoder.scala 71:46]
  wire  func6_op_10000; // @[InstDecoder.scala 72:46]
  wire [4:0] _T_63; // @[InstDecoder.scala 85:33]
  wire  inst_I; // @[InstDecoder.scala 91:39]
  wire  inst_R; // @[InstDecoder.scala 92:39]
  wire  inst_IW; // @[InstDecoder.scala 93:39]
  wire  inst_RW; // @[InstDecoder.scala 94:39]
  wire  _T_94; // @[InstDecoder.scala 49:40]
  wire  _T_98; // @[InstDecoder.scala 46:25]
  wire  _T_100; // @[InstDecoder.scala 46:25]
  wire  _T_102; // @[InstDecoder.scala 46:25]
  wire  _T_104; // @[InstDecoder.scala 46:25]
  wire  _T_106; // @[InstDecoder.scala 46:25]
  wire  _T_112; // @[InstDecoder.scala 46:25]
  wire  _T_114; // @[InstDecoder.scala 46:25]
  wire  inst_SLTI; // @[InstDecoder.scala 46:15]
  wire  inst_SLTIU; // @[InstDecoder.scala 46:15]
  wire  inst_XORI; // @[InstDecoder.scala 46:15]
  wire  inst_ORI; // @[InstDecoder.scala 46:15]
  wire  inst_ANDI; // @[InstDecoder.scala 46:15]
  wire  _T_144; // @[InstDecoder.scala 52:15]
  wire  inst_SLLI; // @[InstDecoder.scala 52:44]
  wire  _T_147; // @[InstDecoder.scala 52:15]
  wire  inst_SRLI; // @[InstDecoder.scala 52:44]
  wire  inst_SRAI; // @[InstDecoder.scala 52:44]
  wire  _T_153; // @[InstDecoder.scala 52:15]
  wire  _T_159; // @[InstDecoder.scala 52:15]
  wire  inst_SLL; // @[InstDecoder.scala 52:44]
  wire  _T_162; // @[InstDecoder.scala 52:15]
  wire  inst_SLT; // @[InstDecoder.scala 52:44]
  wire  _T_165; // @[InstDecoder.scala 52:15]
  wire  inst_SLTU; // @[InstDecoder.scala 52:44]
  wire  _T_168; // @[InstDecoder.scala 52:15]
  wire  inst_XOR; // @[InstDecoder.scala 52:44]
  wire  _T_171; // @[InstDecoder.scala 52:15]
  wire  inst_SRL; // @[InstDecoder.scala 52:44]
  wire  inst_SRA; // @[InstDecoder.scala 52:44]
  wire  _T_177; // @[InstDecoder.scala 52:15]
  wire  inst_OR; // @[InstDecoder.scala 52:44]
  wire  _T_180; // @[InstDecoder.scala 52:15]
  wire  inst_AND; // @[InstDecoder.scala 52:44]
  wire  inst_ADDIW; // @[InstDecoder.scala 46:15]
  wire  _T_185; // @[InstDecoder.scala 52:15]
  wire  inst_SLLIW; // @[InstDecoder.scala 52:44]
  wire  _T_188; // @[InstDecoder.scala 52:15]
  wire  inst_SRLIW; // @[InstDecoder.scala 52:44]
  wire  inst_SRAIW; // @[InstDecoder.scala 52:44]
  wire  _T_194; // @[InstDecoder.scala 52:15]
  wire  inst_ADDW; // @[InstDecoder.scala 52:44]
  wire  _T_200; // @[InstDecoder.scala 52:15]
  wire  inst_SLLW; // @[InstDecoder.scala 52:44]
  wire  _T_203; // @[InstDecoder.scala 52:15]
  wire  inst_SRLW; // @[InstDecoder.scala 52:44]
  wire  inst_SRAW; // @[InstDecoder.scala 52:44]
  OneHotDecoder_1 decoder_3_8 ( // @[InstDecoder.scala 41:27]
    .io_in(decoder_3_8_io_in),
    .io_out(decoder_3_8_io_out)
  );
  OneHotEncoder alu_op_encoder ( // @[InstDecoder.scala 288:30]
    .io_in_1(alu_op_encoder_io_in_1),
    .io_in_2(alu_op_encoder_io_in_2),
    .io_in_3(alu_op_encoder_io_in_3),
    .io_in_4(alu_op_encoder_io_in_4),
    .io_in_5(alu_op_encoder_io_in_5),
    .io_in_6(alu_op_encoder_io_in_6),
    .io_in_7(alu_op_encoder_io_in_7),
    .io_in_8(alu_op_encoder_io_in_8),
    .io_in_9(alu_op_encoder_io_in_9),
    .io_in_10(alu_op_encoder_io_in_10),
    .io_in_11(alu_op_encoder_io_in_11),
    .io_in_12(alu_op_encoder_io_in_12),
    .io_in_13(alu_op_encoder_io_in_13),
    .io_in_14(alu_op_encoder_io_in_14),
    .io_out(alu_op_encoder_io_out)
  );
  assign _T_37 = io_inst[31:25]; // @[InstDecoder.scala 69:38]
  assign func7_op_0 = _T_37 == 7'h0; // @[InstDecoder.scala 69:46]
  assign func7_op_100000 = _T_37 == 7'h20; // @[InstDecoder.scala 70:46]
  assign _T_41 = io_inst[31:26]; // @[InstDecoder.scala 71:38]
  assign func6_op_0 = _T_41 == 6'h0; // @[InstDecoder.scala 71:46]
  assign func6_op_10000 = _T_41 == 6'h10; // @[InstDecoder.scala 72:46]
  assign _T_63 = io_inst[6:2]; // @[InstDecoder.scala 85:33]
  assign inst_I = _T_63 == 5'h4; // @[InstDecoder.scala 91:39]
  assign inst_R = _T_63 == 5'hc; // @[InstDecoder.scala 92:39]
  assign inst_IW = _T_63 == 5'h6; // @[InstDecoder.scala 93:39]
  assign inst_RW = _T_63 == 5'he; // @[InstDecoder.scala 94:39]
  assign _T_94 = decoder_3_8_io_out[0]; // @[InstDecoder.scala 49:40]
  assign _T_98 = decoder_3_8_io_out[1]; // @[InstDecoder.scala 46:25]
  assign _T_100 = decoder_3_8_io_out[4]; // @[InstDecoder.scala 46:25]
  assign _T_102 = decoder_3_8_io_out[5]; // @[InstDecoder.scala 46:25]
  assign _T_104 = decoder_3_8_io_out[6]; // @[InstDecoder.scala 46:25]
  assign _T_106 = decoder_3_8_io_out[7]; // @[InstDecoder.scala 46:25]
  assign _T_112 = decoder_3_8_io_out[2]; // @[InstDecoder.scala 46:25]
  assign _T_114 = decoder_3_8_io_out[3]; // @[InstDecoder.scala 46:25]
  assign inst_SLTI = inst_I & _T_112; // @[InstDecoder.scala 46:15]
  assign inst_SLTIU = inst_I & _T_114; // @[InstDecoder.scala 46:15]
  assign inst_XORI = inst_I & _T_100; // @[InstDecoder.scala 46:15]
  assign inst_ORI = inst_I & _T_104; // @[InstDecoder.scala 46:15]
  assign inst_ANDI = inst_I & _T_106; // @[InstDecoder.scala 46:15]
  assign _T_144 = inst_I & _T_98; // @[InstDecoder.scala 52:15]
  assign inst_SLLI = _T_144 & func6_op_0; // @[InstDecoder.scala 52:44]
  assign _T_147 = inst_I & _T_102; // @[InstDecoder.scala 52:15]
  assign inst_SRLI = _T_147 & func6_op_0; // @[InstDecoder.scala 52:44]
  assign inst_SRAI = _T_147 & func6_op_10000; // @[InstDecoder.scala 52:44]
  assign _T_153 = inst_R & _T_94; // @[InstDecoder.scala 52:15]
  assign _T_159 = inst_R & _T_98; // @[InstDecoder.scala 52:15]
  assign inst_SLL = _T_159 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_162 = inst_R & _T_112; // @[InstDecoder.scala 52:15]
  assign inst_SLT = _T_162 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_165 = inst_R & _T_114; // @[InstDecoder.scala 52:15]
  assign inst_SLTU = _T_165 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_168 = inst_R & _T_100; // @[InstDecoder.scala 52:15]
  assign inst_XOR = _T_168 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_171 = inst_R & _T_102; // @[InstDecoder.scala 52:15]
  assign inst_SRL = _T_171 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign inst_SRA = _T_171 & func7_op_100000; // @[InstDecoder.scala 52:44]
  assign _T_177 = inst_R & _T_104; // @[InstDecoder.scala 52:15]
  assign inst_OR = _T_177 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_180 = inst_R & _T_106; // @[InstDecoder.scala 52:15]
  assign inst_AND = _T_180 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign inst_ADDIW = inst_IW & _T_94; // @[InstDecoder.scala 46:15]
  assign _T_185 = inst_IW & _T_98; // @[InstDecoder.scala 52:15]
  assign inst_SLLIW = _T_185 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_188 = inst_IW & _T_102; // @[InstDecoder.scala 52:15]
  assign inst_SRLIW = _T_188 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign inst_SRAIW = _T_188 & func7_op_100000; // @[InstDecoder.scala 52:44]
  assign _T_194 = inst_RW & _T_94; // @[InstDecoder.scala 52:15]
  assign inst_ADDW = _T_194 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_200 = inst_RW & _T_98; // @[InstDecoder.scala 52:15]
  assign inst_SLLW = _T_200 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign _T_203 = inst_RW & _T_102; // @[InstDecoder.scala 52:15]
  assign inst_SRLW = _T_203 & func7_op_0; // @[InstDecoder.scala 52:44]
  assign inst_SRAW = _T_203 & func7_op_100000; // @[InstDecoder.scala 52:44]
  assign io_aluOPCode = alu_op_encoder_io_out; // @[InstDecoder.scala 290:16]
  assign io_regInfos_0_regIdx = io_inst[19:15]; // @[InstDecoder.scala 27:27]
  assign io_regInfos_0_need = 1'h1; // @[InstDecoder.scala 32:25]
  assign io_regInfos_1_regIdx = io_inst[24:20]; // @[InstDecoder.scala 28:27]
  assign io_regInfos_1_need = 1'h1; // @[InstDecoder.scala 33:25]
  assign io_regInfos_2_regIdx = io_inst[31:27]; // @[InstDecoder.scala 29:27]
  assign io_regInfos_2_need = 1'h1; // @[InstDecoder.scala 34:25]
  assign io_regInfos_3_regIdx = io_inst[11:7]; // @[InstDecoder.scala 30:27]
  assign io_regInfos_3_need = 1'h1; // @[InstDecoder.scala 35:25]
  assign decoder_3_8_io_in = io_inst[14:12]; // @[InstDecoder.scala 42:21]
  assign alu_op_encoder_io_in_1 = _T_153 & func7_op_100000; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_2 = inst_SLTI | inst_SLT; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_3 = inst_SLTIU | inst_SLTU; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_4 = inst_XORI | inst_XOR; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_5 = inst_ORI | inst_OR; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_6 = inst_ANDI | inst_AND; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_7 = inst_SLLI | inst_SLL; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_8 = inst_SRLI | inst_SRL; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_9 = inst_SRAI | inst_SRA; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_10 = inst_ADDIW | inst_ADDW; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_11 = _T_194 & func7_op_100000; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_12 = inst_SLLIW | inst_SLLW; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_13 = inst_SRLIW | inst_SRLW; // @[InstDecoder.scala 289:24]
  assign alu_op_encoder_io_in_14 = inst_SRAIW | inst_SRAW; // @[InstDecoder.scala 289:24]
endmodule
